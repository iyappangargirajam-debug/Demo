Checking if Git is working !!
